// Code your design here
module norgate(input a,b, output c);
nor(c,a,b);
endmodule
