//module declaration with IO ports
module nor_gate(input a, b, output y);

//Logic
nor (y,a,b);

//end of the module
endmodule
