// Code your design here
module nandgate(input a,b, output c);
nand(c,a,b);
endmodule
