//module declaration with IO ports
module nand_gate(input a, b, output y);

//Logic
nand (y,a,b);

//end of the module
endmodule
