//module declaration with IO ports
module xor_gate(input a, b, output y);

//Logic
 xor (y,a,b);

//end of the module
endmodule
