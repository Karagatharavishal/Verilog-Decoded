//module declaration with IO ports
module not_gate(input a, output b);

//logic declaration
  not a1(b, a);
endmodule
