// Code your design here
module xorgate(input a,b, output c);
xor(c,a,b);
endmodule
