//module declaration with IO ports
module and_gate(input a, b, output y);

//Logic
and (y,a,b);

//end of the module
endmodule
