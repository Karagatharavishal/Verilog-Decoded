// Code your design here
//module declaration with IO ports
module xnor_gate(input a, b, output y);

//Logic
 xnor (y,a,b);

//end of the module
endmodule
