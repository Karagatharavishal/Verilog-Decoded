//module declaration with IO ports
module or_gate(input a, b, output c);

//logic declaration
  or a1(c,a,b);
endmodule
