module and_gate (input a, b, output y);
and (y,a,b);
endmodule
