// Code your design here
module xnorgate(input a,b, output c);
xnor(c,a,b);
endmodule
